library verilog;
use verilog.vl_types.all;
entity mux_n_to_8_vlg_vec_tst is
end mux_n_to_8_vlg_vec_tst;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY LCD IS
	GENERIC(
		ULTRA_NUMBER : INTEGER := 3;
		CLK_PERIOD_NS : POSITIVE := 20
	);
	PORT(
		CLK : IN STD_LOGIC;
		RST : IN STD_LOGIC;
		COUNT_IN : IN STD_LOGIC_VECTOR(ULTRA_NUMBER * 8 - 1 DOWNTO 0);
		LCD_E  : OUT STD_LOGIC;
		LCD_RS : OUT STD_LOGIC;
		LCD_RW : OUT STD_LOGIC;
		LCD_DB : OUT STD_LOGIC_VECTOR(7 DOWNTO 4)
	);
END ENTITY LCD;

ARCHITECTURE BEHAVIOR OF LCD IS
	-- LCD PART 
	SIGNAL LINE1 : STD_LOGIC_VECTOR(127 DOWNTO 0);
	SIGNAL LINE2 : STD_LOGIC_VECTOR(127 DOWNTO 0);
	SIGNAL LINE1_BUFFER : STD_LOGIC_VECTOR(127 DOWNTO 0);
	SIGNAL LINE2_BUFFER : STD_LOGIC_VECTOR(127 DOWNTO 0);
	SIGNAL ONE_HZ_CLK : STD_LOGIC;
	-- THIS PART
	SIGNAL COUNT_COUNTER_0 : INTEGER RANGE 0 TO 10 := 0;
	SIGNAL COUNT_COUNTER_1 : INTEGER RANGE 0 TO 10 := 0;
	SIGNAL COUNT_COUNTER_2 : INTEGER RANGE 0 TO 10 := 0;

BEGIN
	LCD : ENTITY WORK.LCD16X2_CTRL
     GENERIC MAP (
      CLK_PERIOD_NS => CLK_PERIOD_NS)
     PORT MAP (
      CLK          => CLK,
      RST          => RST,
      LCD_E        => LCD_E,
      LCD_RS       => LCD_RS,
      LCD_RW       => LCD_RW,
      LCD_DB       => LCD_DB,
      LINE1_BUFFER => LINE1_BUFFER,
      LINE2_BUFFER => LINE2_BUFFER);
		
	DIVIDER : ENTITY WORK.FREQUENCY_DIVIDER
     PORT MAP (
		  CLK        => CLK,				-- CLOCK FROM OSCILLATOR
		  ONE_HZ_CLK => ONE_HZ_CLK);	-- 1 HZ CLOCK
		  
	LINE1(127 DOWNTO 120) <= X"4D"; 
   LINE1(119 DOWNTO 112) <= X"49";
   LINE1(111 DOWNTO 104) <= X"4E";  
   LINE1(103 DOWNTO 96)  <= X"49";  
   LINE1(95 DOWNTO 88)   <= X"50";  
   LINE1(87 DOWNTO 80)   <= X"52";  
   LINE1(79 DOWNTO 72)   <= X"4F";  
   LINE1(71 DOWNTO 64)   <= X"4A";
   LINE1(63 DOWNTO 56)   <= X"2E";  
   LINE1(55 DOWNTO 48)   <= X"20";  
   LINE1(47 DOWNTO 40)   <= X"48";  
   LINE1(39 DOWNTO 32)   <= X"49";  
   LINE1(31 DOWNTO 24)   <= X"47";  
   LINE1(23 DOWNTO 16)   <= X"48";  
   LINE1(15 DOWNTO 8)    <= X"4C";
   LINE1(7 DOWNTO 0)     <= X"56";
		  
	PROCESS(ONE_HZ_CLK)
	BEGIN
		IF RISING_EDGE(ONE_HZ_CLK) THEN
			COUNT_COUNTER_0 <= 0;
			COUNT_COUNTER_1 <= 0;
			COUNT_COUNTER_2 <= 0;
			FOR I IN 0 TO ULTRA_NUMBER-1 LOOP
				IF COUNT_IN((I+1)*8-1 DOWNTO I) > X"FF" THEN
					COUNT_COUNTER_0 <= COUNT_COUNTER_0 + 1;
					IF COUNT_COUNTER_0 = 10 THEN
						COUNT_COUNTER_1 <= COUNT_COUNTER_1 + 1;
						COUNT_COUNTER_0 <= 0;
					END IF;
					IF COUNT_COUNTER_1 = 10 THEN
						COUNT_COUNTER_2 <= COUNT_COUNTER_2 + 1;
						COUNT_COUNTER_1 <= 0;
					END IF;
					IF COUNT_COUNTER_2 = 10 THEN
						COUNT_COUNTER_0 <= 0;
						COUNT_COUNTER_1 <= 0;
						COUNT_COUNTER_2 <= 0;
					END IF;
				END IF;
			END LOOP;
			
			LINE2(127 DOWNTO 120) <= X"4E";
			LINE2(119 DOWNTO 112) <= X"55";
			LINE2(111 DOWNTO 104) <= X"4D";
			LINE2(103 DOWNTO 96)  <= X"42";
			LINE2(95 DOWNTO 88)   <= X"45";
			LINE2(87 DOWNTO 80)   <= X"52";
			LINE2(79 DOWNTO 72)   <= X"20";
			LINE2(71 DOWNTO 64)   <= X"55";
			LINE2(63 DOWNTO 56)   <= X"4C";
			LINE2(55 DOWNTO 48)   <= X"54";
			LINE2(47 DOWNTO 40)   <= X"20";
			LINE2(39 DOWNTO 32)   <= X"3A";
			LINE2(31 DOWNTO 24)   <= X"20";
			LINE2(23 DOWNTO 16)   <= STD_LOGIC_VECTOR(TO_UNSIGNED(COUNT_COUNTER_2, 8));
			LINE2(15 DOWNTO 8)    <= STD_LOGIC_VECTOR(TO_UNSIGNED(COUNT_COUNTER_1, 8));
			LINE2(7 DOWNTO 0)     <= STD_LOGIC_VECTOR(TO_UNSIGNED(COUNT_COUNTER_0, 8));
		END IF;
	END PROCESS;
	LINE1_BUFFER <= LINE1;
   LINE2_BUFFER <= LINE2;
END ARCHITECTURE BEHAVIOR;